library verilog;
use verilog.vl_types.all;
entity ALU is
    port(
        clk             : in     vl_logic;
        S               : in     vl_logic_vector(7 downto 0);
        AC              : out    vl_logic_vector(39 downto 0);
        MQ              : out    vl_logic_vector(39 downto 0);
        MBR             : out    vl_logic_vector(39 downto 0)
    );
end ALU;
